// Instruction Decoder
module instr_Decoder (
	input[8:0] mach_code,
	
);